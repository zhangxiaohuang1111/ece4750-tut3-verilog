//========================================================================
// RegIncr3stage
//========================================================================
// Three-stage registered incrementer that uses structural composition to
// instantitate and connect two instances of the single-stage registered
// incrementer.

`ifndef TUT3_VERILOG_REGINCR_REG_INCR_3STAGE_V
`define TUT3_VERILOG_REGINCR_REG_INCR_3STAGE_V

`include "tut3_verilog/regincr/RegIncr.v"

module tut3_verilog_regincr_RegIncr3stage
(
  input  logic       clk,
  input  logic       reset,
  input  logic [7:0] in_,
  output logic [7:0] out
);

  // First stage

  logic [7:0] reg_incr_0_out;
  logic [7:0] reg_incr_1_out;


  tut3_verilog_regincr_RegIncr reg_incr_0
  (
    .clk    (clk),
    .reset  (reset),
    .in_    (in_),
    .out    (reg_incr_0_out)
  );

// Second stage

tut3_verilog_regincr_RegIncr reg_incr_1 
( 
  .clk (clk), 
  .reset (reset), 
  .in_ (reg_incr_0_out), 
  .out (reg_incr_1_out) 
);

tut3_verilog_regincr_RegIncr reg_incr_2
( 
  .clk (clk), 
  .reset (reset), 
  .in_ (reg_incr_1_out), 
  .out (out) 
);
  // ''' TUTORIAL TASK '''''''''''''''''''''''''''''''''''''''''''''''''''
  // This model is incomplete. As part of the tutorial you will need to
  // instantiate and connect the second stage of this two-stage
  // registered incrementer here.
  // '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

`endif /* TUT3_VERILOG_REGINCR_REG_INCR_3STAGE_V */

